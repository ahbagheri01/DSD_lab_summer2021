library verilog;
use verilog.vl_types.all;
entity mode11_module_vlg_vec_tst is
end mode11_module_vlg_vec_tst;
