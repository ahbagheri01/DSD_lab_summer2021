library verilog;
use verilog.vl_types.all;
entity recognizer_vlg_check_tst is
    port(
        mode3           : in     vl_logic;
        mode11          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end recognizer_vlg_check_tst;
