library verilog;
use verilog.vl_types.all;
entity mode_vlg_vec_tst is
end mode_vlg_vec_tst;
