library verilog;
use verilog.vl_types.all;
entity waiting_room_vlg_vec_tst is
end waiting_room_vlg_vec_tst;
