library verilog;
use verilog.vl_types.all;
entity onebit_comparator_tb is
end onebit_comparator_tb;
