library verilog;
use verilog.vl_types.all;
entity recognizer_vlg_vec_tst is
end recognizer_vlg_vec_tst;
