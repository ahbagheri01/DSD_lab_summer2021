library verilog;
use verilog.vl_types.all;
entity JK_reset_ff_vlg_vec_tst is
end JK_reset_ff_vlg_vec_tst;
