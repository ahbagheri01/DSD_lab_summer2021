library verilog;
use verilog.vl_types.all;
entity onebit_comprator_tb is
end onebit_comprator_tb;
