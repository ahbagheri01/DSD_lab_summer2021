library verilog;
use verilog.vl_types.all;
entity fourbit_comparator_tb is
end fourbit_comparator_tb;
